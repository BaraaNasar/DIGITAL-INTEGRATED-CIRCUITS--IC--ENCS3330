*** SPICE deck for cell PLatch{sch} from library inv
*** Created on Mon Jan 08, 2024 11:08:13
*** Last revised on Thu Aug 22, 2024 03:00:45
*** Written on Thu Aug 22, 2024 03:00:58 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT inv__inv FROM CELL inv{sch}
.SUBCKT inv__inv in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd NMOS L=0.6U W=3U
Mpmos@0 vdd in out vdd PMOS L=0.6U W=3U
.ENDS inv__inv

.global gnd vdd

*** TOP LEVEL CELL: PLatch{sch}
Mnmos@0 out_1210880 net@3 d gnd NMOS L=0.6U W=3U
Mnmos@1 net@50 clk out_1210880 gnd NMOS L=0.6U W=3U
Mpmos@0 out_1210880 clk d vdd PMOS L=0.6U W=3U
Mpmos@1 net@50 net@3 out_1210880 vdd PMOS L=0.6U W=3U
Xinv@1 out_1210880 net@14 inv__inv
Xinv@2 net@14 net@50 inv__inv
Xinv@3 clk net@3 inv__inv

* Spice Code nodes in cell cell 'PLatch{sch}'
vd clk 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb d 0 DC pwl 30n 0 50n 5 120n 5 130n 0
cload out_1210880 0 200fF
.measure tran c_out v(out_1210880) val=4.5 fall=1 td=2ns trag v(out_1210880) val=0.5 fall=1
.measure tran d_out v(out_1210880) val=0.5 rise=1 td=2ns trag v(out_1210880) val=4.5 rise=1
.tran 200n
.include C:\Users\USER\OneDrive\Documents\C5_models.txt
.END
