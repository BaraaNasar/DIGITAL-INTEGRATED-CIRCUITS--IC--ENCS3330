*** SPICE deck for cell NLatch{sch} from library inv
*** Created on Fri Jan 05, 2024 23:59:42
*** Last revised on Thu Aug 22, 2024 02:34:22
*** Written on Thu Aug 22, 2024 02:49:27 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT inv__inv FROM CELL inv{sch}
.SUBCKT inv__inv in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd NMOS L=0.6U W=3U
Mpmos@0 vdd in out vdd PMOS L=0.6U W=3U
.ENDS inv__inv

.global gnd vdd

*** TOP LEVEL CELL: NLatch{sch}
Mnmos@0 out_1210880 clk d gnd NMOS L=0.6U W=3U
Mnmos@1 net@67 net@45 out_1210880 gnd NMOS L=0.6U W=3U
Mpmos@0 out_1210880 net@45 d vdd PMOS L=0.6U W=3U
Mpmos@1 net@67 clk out_1210880 vdd PMOS L=0.6U W=3U
Xinv@0 clk net@45 inv__inv
Xinv@1 out_1210880 net@49 inv__inv
Xinv@2 net@49 net@67 inv__inv

* Spice Code nodes in cell cell 'NLatch{sch}'
vd clk 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb d 0 DC pwl 30n 0 50n 5 120n 5 130n 0
cload out_1210880 0 200fF
.measure tran c_out v(out_1210880) val=4.5 fall=1 td=2ns trag v(out_1210880) val=0.5 fall=1
.measure tran d_out v(out_1210880) val=0.5 rise=1 td=2ns trag v(out_1210880) val=4.5 rise=1
.tran 200n
.include C:\Users\USER\OneDrive\Documents\C5_models.txt
.END
